module vplt

fn vplt() {}